Ex4_6.CIR Drain-feedback bias
vi 1 0 0V ; Value inconsequential
CC 1 2 100uF ; Value inconsequential
RF 2 3 50MEGohm
RL 3 4 3kohm
VDD 4 0 15V
M 3 2 0 0 NMOSG
.MODEL NMOSG NMOS (Vto=4V Kp=0.0008ApVsq
+ Rd=1ohm Rg=1kohm)
.DC VDD 15V 15V 1V
.PRINT DC ID(M) V(2) V(3)
.PROBE
.END

