Prb5_21.CIR
VCC 2 0 15V
VEE 0 7 4V
VIC 3 4 0V
R1 1 0 100ohm
R2 2 1 20kohm
RC 2 3 15kohm
RE 5 6 200ohm
RD 6 7 2kohm
D 0 6 DMOD
Q 4 1 5 QNPNG
.MODEL DMOD D()
.MODEL QNPNG NPN(Is=10fA Ikf=150mA Isc=10fA Bf=150
+ Br=3 Rb=1ohm Rc=1ohm Va=75V Cjc=10pF Cje=15pF)
.DC TEMP 25 125 5
.PROBE
.END
