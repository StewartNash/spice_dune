Ex9_11.CIR
vs 1 0 SIN(0V 0.5V 1kHz)
R2 2 0 1kohm
R2 3 2 10kohm
XA 1 2 3 0 OPAMP
.SUBCKT OPAMP 1   2    3   4
*       Model Inv NInv Out Com
Rd 1 2 500kohm
E 5 4 (1,2) -1e5
Ro 5 3 100ohm
.ENDS OPAMP
.TRAN 1us 2ms
.PROBE
.END

