Ex4_1a..CIR - JFET drain characteristics
vGS 1 0 0V
vDS 2 0 0V
J 2 1 0 NJFET
.MODEL NJFET NJF ( Vto=-4V Beta=0.0005ApVsq
+ Rd=1ohm Rs=1ohm CGS=2pF CGD=2pF)
.DC vDS 0V 25V 0.5V vGS 0V -4V 0.5V
.PROBE
.END
