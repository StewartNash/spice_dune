Prb10_12.CIR
* BOOST CONVERTERRRR
* D=DUTY CYCLE, fs=SWITCHING FREQUENCY
.PARAM D=0.25 fs=20e3Hz
V1 1 0 DC 15V
SW 2 0 4 0 VCS
VSW 4 0 PULSE(0V 1V 0s 5ns 5ns {D/fs} {1/fs})
L 1 2 50uH IC=1.657A
D 2 3 DMOD
C 3 0 100uF IC=20.05V
RL 3 0 7.5ohm
.MODEL DMOD D(N=0.01)
.MODEL VCS VSWITCH(RON=1e-6ohm)
.TRAN 1us 0.25ms 0s 100ns UIC
.PROBE
.END
