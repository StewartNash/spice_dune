* ex_09_12.cir
VS 1 0 AC 1
R1 1 2 1k
R 2 3 10k
C 2 3 0.1u
XA 2 0 3 0 OPAMP
* ------------------
* Op-amp macro-model
* Ideal op-amp subcircuit
.SUBCKT OPAMP 1 2 3 4
* Pins: 1=Inv, 2=NonInv, 3=Out, 4=Common
Rd 1 2 500k
E1 5 4 1 2 -1e5
Ro 5 3 100
.ENDS OPAMP
* ------------------
.AC DEC 200 10 10k
.control
run
shell mkdir -p plots
set hcopydev=png
hardcopy plots/ex_09_12.png db(v(3)/v(1))
quit
.endc
.end

