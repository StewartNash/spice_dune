Prb10_15.CIR
* BUCK-BOOST CONVERTER
* D=DUTY CYLE, fs=SWITCHING FREQUENCY
.PARAM D=0.4 fs=30e3Hz
V1 1 0 DC 15V
SW 1 2 4 2 VCS
VSW 4 2 PULSE(0V 1V 0S 5ns 5ns {D/fs} {1/fs})
L 2 0 70uH IC=0.229A
D 3 2 DMOD
C 0 3 100uF IC=10.02V
RL 0 3 10ohm
.MODEL DMOD D(N=0.01)
.MODEL VCS VSWITCH(RON=1e-6ohm)
.TRAN 1us 0.166667ms 0s 100ns UIC
.PROBE
.END
