* ex8_9_ngspice.cir
* BJT amplifier AC analysis

VI 1 0 AC 0.25

R1 1 0 1k
R2 1 0 16k

VSEN 1 2 DC 0
RHIE 2 3 200
FHFE 3 4 VSEN 90

RE 3 0 500
CE 3 0 330u

RC 4 0 1k
RL 4 0 10k

.AC DEC 25 10 10k

.control
set filetype=ascii
run

* --- Define vectors explicitly ---
let gain_db = db(v(4)/v(1))
let phase_deg = phase(v(4)/v(1))

* --- Write RAW file (optional but safe) ---
write ex8_9_ac.raw

* --- Export ASCII data ---
wrdata ex8_9_ac.dat frequency gain_db phase_deg

quit
.endc

.end

