Prb6_25.CIR
vs 1 0 SIN(0 10mV 10kHz)
VCC 5 0 DC 1115V
CC1 1 2 100uF
CC2 3 4 100uF
CC3 6 8 100uF
CE 7 0 100uF
R11 2 0 100kohm
R12 5 2 90kohm
R22 5 4 90kohm
R21 4 0 10kohm
RE 3 0 9kohm
RC 5 6 5kohm
RL 8 0 5kohm
RE2 7 0 600ohm
Q1 5 2 3 QNPN
Q2 6 4 7 QNPN
.MODEL QNPN NPN()
.PROBE
.TRAN 5us 0.2ms 0s 1us
.END
