Prb6_20.CIR
vs 1 0 SIN(0V 1V 1kHz)
RE 1 0 3.3kohms
Rhib 1 2 25ohms
Vsen 2 0 DC 0V
Fhfb 3 0 Vsen -0.99
Rhob 3 0 {1/1e-6S}
RC 3 0 2.2kohms
RL 3 0 1.1kohms
.TRAN 5 us 1ms
.PROBE
.END
