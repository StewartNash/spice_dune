Ex10_5.CIR
* BUCK CONVERTER
* D=DUTY CYCLE, fs=SWITCHING FREQUENCY
.PARAM D=-.5 fs=25e3Hz
V1 1 0 DC 12V
SW 1 2 4 2 VCS
VSW 4 2 PULSE(0V 1V 0s 5ns 5ns {D/fs} {1/fs})
L 2 3 100uH IC=0.6A
D 0 2 DMOD
C 3 0 50uF IC=6V
RL 3 0 5ohm
.MODEL DMOD D(N=0.01)
.MODEL VCS VSWITCH (RON=1e-6ohm)
.TRAN 5us 0.2ms 0s 100ns UIC
.PROBE
.END
