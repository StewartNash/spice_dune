Prb2_27.CIR
v 1 0 DC 0V
D1 1 2 DMOD
R1 2 3 6kohm
V1 0 3 DC 5V
D2 1 4 DMOD
R2 4 5 3kohm
V2 5 0 DC 10V
.DC v -10V 25V 0.25V
.MODEL DMOD D ()
.PROBE
.END
