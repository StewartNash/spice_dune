Ex9_12.CIR
vs 1 0 AC 1V
R1 1 2 1kohm
R 2 3 10kohm
C 2 3 0.1uF
XA 2 0 3 0 OPAMP
.SUBCKT OPAMP 1   2    3   4
*       Model Inv NInv Out Com
Rd 1 2 500kohm
E 5 4 (1,2) -1e5
Ro 5 3 100ohm
.ENDS OPAMP
.AC DEC 200 10Hz 10kHz
.PROBE
.END
