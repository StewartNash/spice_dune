Ex5_10.CIR
VBB 0 1 -1.32V
VCC 0 4 -15V
RB 1 2 35kohm
RC 3 4 5kohm
RE 5 0 200ohm
Q 3 2 5 QNPNG
.MODEL QNPNG NPN(Is=10fA Ikf=150mA Isc=10fA Bf=150
+ DEV 50% Br=3 RB=1ohm Rc=1ohm Va=75V Cjc=10pF Cje=15pF)
.DC VCC -15V -15V 1V
.WCASE DC IC(Q) YMAX DEVICES Q
.END
