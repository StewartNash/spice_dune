Prb8_20.CIR
vi 1 0 AC 0.25V
RG 1 0 1Megohm
Cgs 1 0 3pF
Cgd 1 2 2.7pF
Ggm 2 0 (1,0) 0.016
rds 2 0 50kohm
Cds 2 0 1pF
RD 2 0 2kohm
RL 2 0 2kohm
.AC DEC 100 1MegHz 100MegHz
.PROBE
.END
